module Quadratic_Equation ();

endmodule // Quadratic_Equation
